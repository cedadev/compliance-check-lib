netcdf amf_eg_data_1 {
dimensions:
	time = 87 ;
	altitude = 21 ;
	latitude = 1 ;
	longitude = 1 ;
variables:
	double aerosol_backscatter_coefficient(time, altitude) ;
		aerosol_backscatter_coefficient:units = "m-1 sr-1" ;
		aerosol_backscatter_coefficient:long_name = "Attenuated backscatter coefficient" ;
		aerosol_backscatter_coefficient:_FillValue = -1.e+20 ;
		aerosol_backscatter_coefficient:valid_min = 1.e-07 ;
		aerosol_backscatter_coefficient:valid_max = 1. ;
		aerosol_backscatter_coefficient:cell_methods = "time: mean" ;
		aerosol_backscatter_coefficient:coordinates = "latitude longitude" ;
	double altitude(altitude) ;
		altitude:units = "m" ;
		altitude:standard_name = "altitude" ;
		altitude:long_name = "Geometric height above geoid (WGS84)." ;
		altitude:_FillValue = -1.e+20 ;
		altitude:axis = "Z" ;
		altitude:valid_min = 0. ;
		altitude:valid_max = 10263. ;
	int day(time) ;
		day:units = "1" ;
		day:long_name = "Day" ;
		day:valid_min = 1. ;
		day:valid_max = 31. ;
	double day_of_year(time) ;
		day_of_year:units = "1" ;
		day_of_year:long_name = "Day of Year" ;
		day_of_year:valid_min = 1. ;
		day_of_year:valid_max = 366. ;
	int hour(time) ;
		hour:units = "1" ;
		hour:long_name = "Hour" ;
		hour:valid_min = 0. ;
		hour:valid_max = 23. ;
	double latitude(latitude) ;
		latitude:units = "degrees_north" ;
		latitude:standard_name = "latitude" ;
		latitude:long_name = "Latitude" ;
	double longitude(longitude) ;
		longitude:units = "degree_east" ;
		longitude:standard_name = "longitude" ;
		longitude:long_name = "Longitude" ;
	int minute(time) ;
		minute:units = "1" ;
		minute:long_name = "Minute" ;
		minute:valid_min = 0. ;
		minute:valid_max = 59. ;
	int month(time) ;
		month:units = "1" ;
		month:long_name = "Month" ;
		month:valid_min = 1. ;
		month:valid_max = 12. ;
	int qc_flag(time, altitude) ;
		qc_flag:units = "1" ;
		qc_flag:long_name = "Data Quality flag" ;
		qc_flag:valid_min = 1. ;
		qc_flag:valid_max = 3. ;
	double second(time) ;
		second:units = "1" ;
		second:long_name = "Second" ;
		second:valid_min = 0. ;
		second:valid_max = 59.9999 ;
	double time(time) ;
		time:units = "seconds since 1970-01-01 00:00:00 UTC" ;
		time:standard_name = "time" ;
		time:long_name = "Time (seconds since 1970-01-01)" ;
		time:axis = "T" ;
		time:valid_min = 1467331210.67063 ;
		time:valid_max = 1467417595.78003 ;
		time:calendar = "julian" ;
	int year(time) ;
		year:units = "1" ;
		year:long_name = "Year" ;
		year:valid_min = 1900. ;
		year:valid_max = 2100. ;

// global attributes:
		:Conventions = "CF-1.6" ;
		:source = "NCAS 905nm Lidar Ceilometer" ;
		:instrument_manufacturer = "Campbell Scientific" ;
		:instrument_model = "CS 135" ;
		:serial_number = "E1002" ;
		:operational_software = "Campbell Scientific firmware" ;
		:operational_software_version = "No version number" ;
		:creator_name = "B.Brooks" ;
		:creator_email = "barbara.brooks@ncas.ac.uk" ;
		:creator_url = "https://amf.ncas.ac.uk" ;
		:institution = "National Centre for Atmospheric Science (NCAS)" ;
		:processing_level = 2 ;
		:processing_software = "Matlab R2013b using Parse_Ceilometer_v1" ;
		:processing_software_version = "v1" ;
		:calibration_sensitivity = "\"Calibrated to manufacturers standard:0.25%, 4.6 m\"" ;
		:calibration_certification_date = "not known" ;
		:calibration_certification_url = "not applicable" ;
		:sampling_interval = "10 seconds" ;
		:averaging_interval = "10 seconds" ;
		:data_set_version = "1.2" ;
		:data_product_level = "1" ;
		:last_revised_date = "2017-02-25T13:14:16" ;
		:project = "Dynamics-aerosol-chemistry-cloud interactions in West Africa. (DACCIWA)" ;
		:project_principle_investigator = "Peter Knippertz" ;
		:project_principle_investigator_contact = "peter.knippertz@kit.edu" ;
		:licence = "Data usage licence - UK Government Open Licence agreement: http://www.nationalarchives.gov.uk/doc/open-government-licence" ;
		:acknowledgement = "Acknowledgement of NCAS as the data provider is required whenever and wherever this data is used" ;
		:platform_type = "stationary_platform" ;
		:platform_name = "kumasi" ;
		:title = "Profiles of attenuated aerosol backscatter coefficient from the NCAS 905nm Lidar Ceilometer at KNUST, Kumasi, Ghana." ;
		:feature_type = "timeSeriesProfile" ;
		:start_time = "2016-07-01T00:00:10" ;
		:end_time = "2016-07-01T23:59:55" ;
		:platform_location = "06 40 46.6 N (6.67961), 01 33 36.4 W (-1.56011)" ;
		:platform_height = "263m" ;
		:location_keywords = "africa, ghana, kumasi, knust" ;
		:history = "Thu Dec  7 00:21:17 2017: ncks -d time,,,100 -d altitude,,,100 orig/ncas-ceil-1_kumasi_20160701_backscatter_v1.2.nc ncas-ceil-1_kumasi_20160701_backscatter_v1.2.nc\n",
			"Data collected June - July 2016, processed & QC\'d Oct 2016. v1.1 minor revision to correct Cf compliance issues. V1.2 corrects for time unit error." ;
		:comment = "" ;
		:qc_flag_comment = "integer in the range 0 - 3" ;
		:qc_flag_value_0_description = "not used" ;
		:qc_flag_value_1_description = "good data" ;
		:qc_flag_value_1_assessment = "good data" ;
		:qc_flag_value_2_description = "Attenuated aerosol backscatter coefficient outside instrument operational range" ;
		:qc_flag_value_2_assessment = "bad data" ;
		:qc_flag_value_3_description = "Time stamp error" ;
		:qc_flag_value_3_assessment = "suspect data" ;
		:NCO = "\"4.5.5\"" ;
data:

 aerosol_backscatter_coefficient =
  0.0524286, 0.000194, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.0524286, _, 2.09e-05, _, _, _, _, _, _, 0.0008444, _, _, 0.004125, _, _, 
    _, _, _, _, _, 0.0097765,
  0.0524286, 0.0001657, 6.05e-05, 2.24e-05, 1.42e-05, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.0524286, 7.38e-05, 6.26e-05, _, _, _, 5.66e-05, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.0524286, 2.9e-05, 4.85e-05, _, _, _, _, _, _, _, 0.0014832, _, _, _, _, 
    _, _, _, _, _, _,
  0.0524286, 3.74e-05, _, _, _, 0.0004903, _, _, _, _, _, 0.0005795, 
    0.0033188, 0.0004822, _, _, _, _, _, _, _,
  0.0524286, 3.75e-05, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.0524286, 0.0070792, 4.8e-06, 6.8e-05, 6.24e-05, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, 0.0020478, _, _,
  0.0524286, 3.76e-05, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.0524286, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.0524286, 2.96e-05, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.0524286, _, _, 0.000272, _, _, _, _, _, _, _, 0.0018178, _, 0.0010223, 
    0.0084021, _, _, 0.0031374, 0.0076997, 0.0123574, _,
  0.0524286, 6.4e-06, _, _, _, _, _, _, _, _, _, _, _, _, _, 0.0051881, _, _, 
    _, _, _,
  0.0524286, _, _, 0.0001793, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    0.0023437,
  0.0524286, 0.0011493, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.0524286, 0.000553, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.0524286, 0.0002303, 8.36e-05, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0.0524286, _, _, _, _, _, _, _, _, _, 0.0005369, _, _, _, _, _, _, _, _, _, _,
  0.0524286, 2.42e-05, 0.000113, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.0524286, 0.0001706, 6.95e-05, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0.0524286, 4.45e-05, 3.75e-05, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.0524286, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0.0031748, _, _, _,
  0.0524286, _, 0.0002557, 0.000853, _, _, _, _, _, _, _, _, 0.0102515, 
    0.0033534, 0.0047981, 0.0100562, _, _, _, _, 0.0065716,
  0.0524286, 0.000126, _, _, _, 0.0005642, _, _, 0.0128539, _, _, 0.0130277, 
    0.0204511, _, _, _, 0.0345565, _, _, _, _,
  0.0524286, 0.0002992, _, _, _, _, _, 0.0028505, _, _, _, _, 0.0074042, _, 
    _, _, 0.0030545, _, _, _, _,
  0.0524286, 0.000101, _, _, _, _, 0.0005933, _, 0.0038038, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.0524286, 8.48e-05, _, 4.04e-05, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.0524286, 0.0001514, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.0524286, 0.0001611, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.0524286, 0.0005772, _, 0.0016133, _, 0.0010251, _, 0.0041545, _, _, _, _, 
    _, _, _, 0.0024391, _, 0.0496265, _, _, _,
  0.0524286, 4.35e-05, _, _, _, _, _, _, _, _, _, _, _, _, _, 0.0074851, _, 
    0.0339517, _, _, 0.0096563,
  0.0524286, 0.000623, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.0524286, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.0524286, 0.0005255, _, _, 0.0090603, _, _, 0.004182, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.0524286, _, _, 0.0003082, _, _, _, _, _, 0.0109324, _, _, _, _, _, _, _, 
    _, _, _, _,
  0.0524286, _, _, _, 0.0043204, _, 0.0047436, _, _, _, 0.0063895, _, _, _, 
    _, _, _, _, _, _, _,
  0.0524286, 0.0003729, _, _, _, _, _, _, _, _, _, _, 0.0109566, _, _, _, _, 
    0.0203859, _, _, _,
  0.0524286, 0.0444614, 0.0004248, _, _, _, 0.0056015, 0.005767, _, _, _, _, 
    _, _, _, _, _, _, 0.0048523, _, _,
  0.0524286, 0.0246982, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.0524286, _, _, _, _, _, _, _, _, 0.0043347, _, _, 0.0020543, _, _, _, 
    0.0140843, _, _, _, _,
  0.0524286, 0.0003715, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    0.0163957, 0.0524286, _, _,
  0.0524286, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.0524286, _, _, _, 0.0005035, _, 0.0009759, 0.0023198, _, _, _, _, _, _, 
    _, _, _, 0.0143659, 0.0078304, _, _,
  0.0524286, 9.58e-05, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.0524286, _, _, _, _, _, _, 0.0026811, _, _, _, _, 0.01029, _, _, _, _, _, 
    _, _, _,
  0.0524286, _, _, _, _, _, _, 0.0012192, _, 0.0042093, _, _, _, _, _, 
    0.0078678, _, _, _, _, _,
  0.0524286, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.0524286, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.0524286, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.0524286, _, 0.0001086, _, _, _, _, _, _, 0.0013804, _, _, 0.0070838, _, 
    _, _, _, _, _, _, _,
  0.0524286, 4.96e-05, _, _, _, _, _, 0.0048612, _, _, _, 0.0024862, _, 
    0.0046182, _, _, 0.004115, _, _, 0.0216256, _,
  0.0524286, 3.24e-05, 0.0003468, _, _, _, _, _, 0.0012044, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.0524286, 1.68e-05, _, _, _, 0.0056445, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0.0524286, 9.6e-06, _, _, _, _, _, 0.0002567, _, _, _, _, 0.0006097, _, _, 
    _, _, _, _, _, _,
  0.0524286, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0.0071724, _, _,
  0.0524286, 2.2e-05, _, 0.0002495, 0.000581, _, _, 0.0044658, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.0524286, 9.77e-05, _, _, _, _, _, _, _, _, _, _, _, _, _, 0.007564, _, 
    0.0055848, _, _, _,
  0.0524286, 0.0001103, _, _, _, _, _, _, _, _, _, _, 0.0021624, _, _, _, 
    0.0051659, 0.0042367, _, _, _,
  0.0524286, 0.0001023, _, _, _, _, _, _, _, _, 0.0018755, _, _, 0.0008484, 
    _, 0.006364, _, _, _, _, _,
  0.0524286, 0.0001059, _, 7.29e-05, _, _, _, _, _, _, _, _, _, _, _, _, 
    0.002576, 0.0008485, _, _, _,
  0.0524286, 0.000102, _, _, _, _, _, _, _, _, _, _, _, _, _, 0.0028061, _, 
    _, _, _, _,
  0.0524286, 9.04e-05, _, _, 0.000637, _, 0.0007833, 0.0005713, 0.0002929, _, 
    _, _, 0.0038884, _, _, _, 0.0113602, _, _, _, _,
  0.0524286, 8.41e-05, _, _, 0.0001457, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0.0524286, 5.09e-05, _, _, _, _, _, _, _, 0.0003589, _, _, _, _, _, _, _, 
    _, _, _, _,
  0.0524286, 7.46e-05, _, _, _, 0.0034143, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0.0524286, 6.42e-05, 1.75e-05, _, _, _, _, _, _, 0.0001112, _, _, _, _, _, 
    _, _, 0.0045945, 0.0004295, _, _,
  0.0524286, 0.0001106, 8.85e-05, _, 2.05e-05, 3.14e-05, _, _, _, 0.0008429, 
    _, 0.0013465, _, _, _, _, _, 0.0029625, _, _, _,
  0.0524286, 7.4e-05, 4.18e-05, 1.61e-05, _, _, 0.0001854, _, _, _, _, _, 
    8.2e-05, _, 0.0001879, _, _, _, _, _, _,
  0.0524286, 7.14e-05, 5.12e-05, 2.2e-05, 7.35e-05, _, _, _, _, 0.0004177, _, 
    0.0004921, _, _, _, 0.0009084, _, _, _, 0.0008655, _,
  0.0524286, 7.01e-05, 5.16e-05, 5e-05, 2.11e-05, _, _, _, 5.51e-05, _, _, 
    4.78e-05, _, _, _, _, _, _, _, _, _,
  0.0524286, 5.58e-05, 6.5e-05, _, _, _, _, 0.000351, _, 8.63e-05, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.0524286, 4.7e-05, 4.4e-05, 3.37e-05, _, _, _, _, _, _, _, _, _, _, 
    7.46e-05, _, _, _, _, _, _,
  0.0524286, 7.07e-05, 5.15e-05, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    0.0002236, _, _, _,
  0.0524286, 5.24e-05, 5.97e-05, 5.39e-05, _, _, _, _, _, _, _, 0.0001625, _, 
    _, _, _, _, _, 0.0001259, _, _,
  0.0524286, 0.0001321, 4.71e-05, 5.23e-05, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.0524286, 6.09e-05, 4.86e-05, _, 1.24e-05, _, _, _, 5.24e-05, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.0524286, 6.54e-05, 5.53e-05, 1.17e-05, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.0524286, 8.31e-05, 6.2e-05, _, _, _, _, _, _, _, _, _, _, _, 0.0002598, 
    _, _, _, _, _, _,
  0.0524286, 8.77e-05, 4.66e-05, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.0524286, 0.0001001, 5.79e-05, 6.36e-05, _, _, _, _, _, _, _, _, _, _, 
    8.14e-05, _, _, _, _, _, _,
  0.0524286, 8.26e-05, 6.21e-05, 5.29e-05, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.0524286, 0.0001127, 7.54e-05, _, _, _, _, _, _, _, _, _, 8.99e-05, _, _, 
    _, _, _, 0.0005286, _, _,
  0.0524286, 0.0001112, 6.72e-05, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0.0524286, 0.0098896, 5.64e-05, _, 0.0001116, _, _, _, 0.0002174, _, _, _, 
    _, 0.0003792, _, _, _, _, 0.0001567, _, _,
  0.0524286, 0.000177, 7.37e-05, 2.86e-05, 5.52e-05, _, _, _, _, _, 
    0.0001024, _, _, _, _, 0.0002552, _, _, _, _, _,
  0.0524286, 0.000398, 6.93e-05, _, 7.4e-06, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, 0.000207, _,
  0.0524286, 0.0001126, 4.5e-05, _, _, _, 5.03e-05, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _ ;

 altitude = 265.5, 765.5, 1265.5, 1765.5, 2265.5, 2765.5, 3265.5, 3765.5, 
    4265.5, 4765.5, 5265.5, 5765.5, 6265.5, 6765.5, 7265.5, 7765.5, 8265.5, 
    8765.5, 9265.5, 9765.5, 10265.5 ;

 day = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 day_of_year = 183.000123502687, 183.011694011046, 183.023267395096, 
    183.034839822561, 183.046528865001, 183.058100031922, 183.069670370547, 
    183.081243609311, 183.092815204524, 183.10438588378, 183.115959245828, 
    183.127532846062, 183.139102185378, 183.150674283504, 183.162250009016, 
    183.173819859279, 183.185390525497, 183.196963115362, 183.208535791025, 
    183.220106619643, 183.231678684708, 183.243250679108, 183.254825281445, 
    183.266398713225, 183.277969841147, 183.289539205725, 183.301114186412, 
    183.312683661468, 183.324255404761, 183.335827549105, 183.347402114305, 
    183.358971632901, 183.37054832885, 183.38211682823, 183.393687817501, 
    183.405260321451, 183.416831928655, 183.42840469908, 183.439977839123, 
    183.451550909784, 183.463120228727, 183.474693319993, 183.486264379928, 
    183.497839554679, 183.509410108789, 183.520982373157, 183.532556238468, 
    183.544124859734, 183.555698163575, 183.567270514555, 183.578841057839, 
    183.590413870057, 183.601986348978, 183.613560447586, 183.625129484804, 
    183.636701517738, 183.648274182342, 183.659845750197, 183.671535674832, 
    183.683106088545, 183.694680573768, 183.706252141623, 183.717937541194, 
    183.729509577621, 183.741082462715, 183.752653758391, 183.764228152111, 
    183.775801519281, 183.787369976053, 183.798941944027, 183.810522233602, 
    183.822087632143, 183.833660762408, 183.845230378909, 183.856803539558, 
    183.868377562496, 183.879946806584, 183.891518930322, 183.903090997483, 
    183.91466312937, 183.926235251944, 183.937807378941, 183.949379725382, 
    183.96095323097, 183.972525038291, 183.984095712309, 183.995667788084 ;

 hour = 0, 0, 0, 0, 1, 1, 1, 1, 2, 2, 2, 3, 3, 3, 3, 4, 4, 4, 5, 5, 5, 5, 6, 
    6, 6, 6, 7, 7, 7, 8, 8, 8, 8, 9, 9, 9, 10, 10, 10, 10, 11, 11, 11, 11, 
    12, 12, 12, 13, 13, 13, 13, 14, 14, 14, 15, 15, 15, 15, 16, 16, 16, 16, 
    17, 17, 17, 18, 18, 18, 18, 19, 19, 19, 20, 20, 20, 20, 21, 21, 21, 21, 
    22, 22, 22, 23, 23, 23, 23 ;

 latitude = 6.67961 ;

 longitude = -1.56011 ;

 minute = 0, 16, 33, 50, 7, 23, 40, 56, 13, 30, 46, 3, 20, 36, 53, 10, 26, 
    43, 0, 16, 33, 50, 6, 23, 40, 56, 13, 30, 46, 3, 20, 36, 53, 10, 26, 43, 
    0, 16, 33, 50, 6, 23, 40, 56, 13, 30, 46, 3, 20, 36, 53, 10, 26, 43, 0, 
    16, 33, 50, 7, 23, 40, 57, 13, 30, 47, 3, 20, 37, 53, 10, 27, 43, 0, 17, 
    33, 50, 7, 23, 40, 57, 13, 30, 47, 3, 20, 37, 53 ;

 month = 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 
    7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 
    7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 
    7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7 ;

 qc_flag =
  1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 2, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 2, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 2, 2, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 2, 2, 2, 1, 2, 2, 2, 2, 2, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 2, 2, 2, 2, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 2, 2, 2, 2, 2, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 2, 2, 2, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 ;

 second = 10.670629, 50.362555, 30.302938, 10.160667, 0.093937, 39.842757, 
    19.520012, 59.447843, 39.233674, 18.940357, 58.878837, 38.837897, 
    18.428817, 58.258094, 38.400782, 18.035842, 57.741407, 37.613167, 
    17.492348, 57.211941, 37.038357, 16.858675, 56.904319, 36.848826, 
    16.594275, 56.187377, 36.265706, 15.868352, 55.666976, 35.500247, 
    15.542678, 55.14908, 35.375611, 14.893955, 54.627433, 34.491778, 
    14.27864, 54.166001, 34.085305, 13.998605, 53.587763, 33.502851, 
    13.242428, 53.337527, 33.033401, 12.877036, 52.859007, 32.387885, 
    12.321335, 52.172457, 31.867395, 11.758373, 51.620556, 31.622675, 
    11.187483, 51.011135, 30.88935, 10.672819, 0.682305, 40.366051, 
    20.401569, 0.185032, 49.803563, 29.627504, 9.524775, 49.28472, 29.312339, 
    9.251265, 48.765935, 28.58396, 9.120979, 48.371416, 28.28987, 7.904741, 
    47.825816, 27.821403, 7.404086, 47.235582, 27.062179, 6.894382, 
    46.725765, 26.557541, 6.408275, 46.359159, 26.163306, 5.869541, 45.696888 ;

 time = 1467331210.67063, 1467332210.36255, 1467333210.30294, 
    1467334210.16067, 1467335220.09394, 1467336219.84276, 1467337219.52002, 
    1467338219.44784, 1467339219.23367, 1467340218.94036, 1467341218.87884, 
    1467342218.8379, 1467343218.42882, 1467344218.25809, 1467345218.40078, 
    1467346218.03584, 1467347217.7414, 1467348217.61317, 1467349217.49234, 
    1467350217.21194, 1467351217.03836, 1467352216.85868, 1467353216.90432, 
    1467354216.84882, 1467355216.59427, 1467356216.18737, 1467357216.26571, 
    1467358215.86835, 1467359215.66697, 1467360215.50024, 1467361215.54268, 
    1467362215.14908, 1467363215.37561, 1467364214.89396, 1467365214.62743, 
    1467366214.49177, 1467367214.27864, 1467368214.166, 1467369214.0853, 
    1467370213.99861, 1467371213.58776, 1467372213.50285, 1467373213.24243, 
    1467374213.33752, 1467375213.0334, 1467376212.87704, 1467377212.859, 
    1467378212.38788, 1467379212.32133, 1467380212.17246, 1467381211.8674, 
    1467382211.75837, 1467383211.62055, 1467384211.62267, 1467385211.18749, 
    1467386211.01113, 1467387210.88935, 1467388210.67282, 1467389220.68231, 
    1467390220.36605, 1467391220.40157, 1467392220.18504, 1467393229.80356, 
    1467394229.62751, 1467395229.52478, 1467396229.28472, 1467397229.31234, 
    1467398229.25127, 1467399228.76593, 1467400228.58396, 1467401229.12098, 
    1467402228.37142, 1467403228.28987, 1467404227.90474, 1467405227.82582, 
    1467406227.8214, 1467407227.40409, 1467408227.23558, 1467409227.06218, 
    1467410226.89438, 1467411226.72577, 1467412226.55754, 1467413226.40827, 
    1467414226.35916, 1467415226.16331, 1467416225.86954, 1467417225.69689 ;

 year = 2016, 2016, 2016, 2016, 2016, 2016, 2016, 2016, 2016, 2016, 2016, 
    2016, 2016, 2016, 2016, 2016, 2016, 2016, 2016, 2016, 2016, 2016, 2016, 
    2016, 2016, 2016, 2016, 2016, 2016, 2016, 2016, 2016, 2016, 2016, 2016, 
    2016, 2016, 2016, 2016, 2016, 2016, 2016, 2016, 2016, 2016, 2016, 2016, 
    2016, 2016, 2016, 2016, 2016, 2016, 2016, 2016, 2016, 2016, 2016, 2016, 
    2016, 2016, 2016, 2016, 2016, 2016, 2016, 2016, 2016, 2016, 2016, 2016, 
    2016, 2016, 2016, 2016, 2016, 2016, 2016, 2016, 2016, 2016, 2016, 2016, 
    2016, 2016, 2016, 2016 ;
}
